`include "dma_transaction_thread00.v"
