`include "dma_transaction_thread02.v"
