//`include "dma_transaction_for_thread02.v"
