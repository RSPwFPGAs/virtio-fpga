`include "dma_transaction_thread01.v"
