`include "dma_transaction_thread03.v"
