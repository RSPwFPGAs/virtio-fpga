`timescale 1ns / 100ps

//`include "axi_vip_0_exdes_generic.sv"
`include "axi_vip_0_passthrough_mst_stimulus.sv"
`include "axi_vip_thread00_passthrough_mst_stimulus.sv"
`include "axi_vip_thread01_passthrough_mst_stimulus.sv"
`include "axi_vip_thread02_passthrough_mst_stimulus.sv"
`include "axi_vip_thread03_passthrough_mst_stimulus.sv"
`include "axi_vip_thread04_passthrough_mst_stimulus.sv"
`include "axi_vip_thread05_passthrough_mst_stimulus.sv"
`include "axi_vip_thread06_passthrough_mst_stimulus.sv"
//`include "axi_vip_0_slv_basic_stimulus.sv"

module test_top ();

reg  PCIE_CLK_N;
reg  PCIE_CLK_P;
wire [7:0] PCIE_RX_N;
wire [7:0] PCIE_RX_P;
wire [7:0] PCIE_TX_N;
wire [7:0] PCIE_TX_P;
reg  PERSTN;
reg  FPGA_SYSCLK_N;
reg  FPGA_SYSCLK_P;
reg  RESET;
wire  UART_RXD_OUT;
wire  UART_TXD_IN;
shell_region_wrapper DUT (
  .pci_express_rxn (PCIE_RX_N),
  .pci_express_rxp (PCIE_RX_P),
  .pci_express_txn (PCIE_TX_N),
  .pci_express_txp (PCIE_TX_P),
  .pcie_perstn (PERSTN),
  .pcie_refclk_clk_n (PCIE_CLK_N),
  .pcie_refclk_clk_p (PCIE_CLK_P)
);

// instantiate vip master
//  axi_vip_0_exdes_generic  generic_tb();
  axi_vip_0_passthrough_mst_stimulus mst_axilite_toCSR();  // for initialization of CSR
  axi_vip_thread00_passthrough_mst_stimulus mst_axifull_toDMA_th00();  // for transaction of DMA
  axi_vip_thread01_passthrough_mst_stimulus mst_axifull_toDMA_th01();  // for transaction of DMA
  axi_vip_thread02_passthrough_mst_stimulus mst_axifull_toDMA_th02();  // for transaction of DMA
  axi_vip_thread03_passthrough_mst_stimulus mst_axifull_toDMA_th03();  // for transaction of DMA
  axi_vip_thread04_passthrough_mst_stimulus mst_axifull_toDMA_th04();  // for transaction of DMA
  axi_vip_thread05_passthrough_mst_stimulus mst_axifull_toDMA_th05();  // for transaction of DMA
  axi_vip_thread06_passthrough_mst_stimulus mst_axifull_toDMA_th06();  // for transaction of DMA
//  axi_vip_0_slv_basic_stimulus slv();
    

//////////////////////////////////
// Inter-thread signals

`define CSR_PATH test_top.DUT.shell_region_i.FIM.FIU.feature_ram.virtio_csr_0.inst
`define TH00_PATH test_top.mst_axifull_toDMA_th00
`define TH01_PATH test_top.mst_axifull_toDMA_th01
`define TH02_PATH test_top.mst_axifull_toDMA_th02
`define TH03_PATH test_top.mst_axifull_toDMA_th03
`define TH04_PATH test_top.mst_axifull_toDMA_th04
`define TH05_PATH test_top.mst_axifull_toDMA_th05
`define TH06_PATH test_top.mst_axifull_toDMA_th06

// inter-thread 0-1 signals
reg queue_notify_pending[3];
// make a record of pending notification
always @(posedge `CSR_PATH.clk) begin
  for (int i = 0; i < 3; i++) begin
    if (`CSR_PATH.csr_rst)
      queue_notify_pending[i] = 1'b0;
    else if (`TH00_PATH.queue_notify_set[i])
      queue_notify_pending[i] = 1'b1;
    else if (`TH01_PATH.queue_notify_clr[i])
      queue_notify_pending[i] = 1'b0;
  end
end

// inter-thread 1-2 signals
reg ring_available_pending[3];
// make a record of pending available rings
always @(posedge `CSR_PATH.clk) begin
  for (int i = 0; i < 3; i++) begin
    if (`CSR_PATH.csr_rst)
      ring_available_pending[i] = 1'b0;
    else if (`TH01_PATH.ring_available_set[i])
      ring_available_pending[i] = 1'b1;
    else if (`TH02_PATH.ring_available_clr[i])
      ring_available_pending[i] = 1'b0;
  end
end

reg [15:0] th01_next_avail_idx[3];
// update next available index
always @(*) begin
  for (int i = 0; i < 3; i++) begin
    th01_next_avail_idx[i] = `TH01_PATH.next_avail_idx[i];
  end
end

//typedef bit [16+128-1:0] desc_q [];
//desc_q desc_queue [$];

// inter-thread 2-345 signals
//bit [16+128-1:0] desc_queue_0 [$] = {};
//bit [16+128-1:0] desc_queue_1 [$] = {};
//bit [16+128-1:0] desc_queue_2 [$] = {};
bit [16+128-1:0] desc_queue[3] [$];  // {desc_idx, desc_entry}

// inter-thread 345-6 signals
//bit [16+32-1:0] ring_used_queue_0 [$] = {};
//bit [16+32-1:0] ring_used_queue_1 [$] = {};
//bit [16+32-1:0] ring_used_queue_2 [$] = {};
bit [16+32-1:0] ring_used_queue[3] [$];  // {desc_idx, desc_chain_len}

//// inter-thread 2-6 signals
//reg ring_used_pending[3];
//// make a record of pending used rings
//always @(posedge `CSR_PATH.clk) begin
//  for (int i = 0; i < 3; i++) begin
//    if (`CSR_PATH.csr_rst)
//      ring_used_pending[i] = 1'b0;
//    else if (`TH02_PATH.ring_used_set[i])
//      ring_used_pending[i] = 1'b1;
//    else if (`TH06_PATH.ring_used_clr[i])
//      ring_used_pending[i] = 1'b0;
//  end
//end
//
//reg [15:0] th02_next_avail_idx[3];
//// update next available index
//always @(*) begin
//  for (int i = 0; i < 3; i++) begin
//    th02_next_avail_idx[i] = `TH02_PATH.next_avail_idx[i];
//  end
//end

// Inter-thread signals
/////////////////////////////////////


always
begin
  PCIE_CLK_N = 1;
  #5.0;
  PCIE_CLK_N = 0;
  #5.0;
end
always
begin
  PCIE_CLK_P = 0;
  #5.0;
  PCIE_CLK_P = 1;
  #5.0;
end

always
begin
  FPGA_SYSCLK_N = 0;
  #2.5;
  FPGA_SYSCLK_N = 1;
  #2.5;
end
always
begin
  FPGA_SYSCLK_P = 1;
  #2.5;
  FPGA_SYSCLK_P = 0;
  #2.5;
end

initial
begin
  $display("[%t] : System Reset(test_top/RESET) Is Asserted...", $realtime);
  RESET = 1;
  #5000;
  $display("[%t] : System Reset(test_top/RESET) Is DeAsserted...", $realtime);
  RESET = 0;
end

initial
begin
  $display("[%t] : System Reset(test_top/PERSTN) Is Asserted...", $realtime);
  PERSTN = 0;
  #100;
  $display("[%t] : System Reset(test_top/PERSTN) Is DeAsserted...", $realtime);
  PERSTN = 1;
end

initial begin
  $display("V: testbench init.");
end

endmodule

