`include "dma_transaction_thread06.v"
