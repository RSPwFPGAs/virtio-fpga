//`include "dma_transaction_for_thread04.v"
