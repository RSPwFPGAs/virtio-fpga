//`include "dma_transaction_for_thread03.v"
