//`include "dma_transaction_for_thread06.v"
