//`include "dma_transaction_thread04.v"
