//`include "dma_transaction_for_thread05.v"
