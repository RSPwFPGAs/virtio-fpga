//`include "dma_transaction_thread05.v"
